library verilog;
use verilog.vl_types.all;
entity ula01_vlg_vec_tst is
end ula01_vlg_vec_tst;
