library verilog;
use verilog.vl_types.all;
entity memory5_vlg_vec_tst is
end memory5_vlg_vec_tst;
