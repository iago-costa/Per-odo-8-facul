library verilog;
use verilog.vl_types.all;
entity ula02_vlg_vec_tst is
end ula02_vlg_vec_tst;
