library verilog;
use verilog.vl_types.all;
entity memory2_vlg_vec_tst is
end memory2_vlg_vec_tst;
