library verilog;
use verilog.vl_types.all;
entity shift_register_vlg_vec_tst is
end shift_register_vlg_vec_tst;
