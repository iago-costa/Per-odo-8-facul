library verilog;
use verilog.vl_types.all;
entity memory2_vlg_check_tst is
    port(
        ssd             : in     vl_logic_vector(6 downto 0);
        sampler_rx      : in     vl_logic
    );
end memory2_vlg_check_tst;
