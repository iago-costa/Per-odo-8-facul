library verilog;
use verilog.vl_types.all;
entity memory3_vlg_vec_tst is
end memory3_vlg_vec_tst;
