library verilog;
use verilog.vl_types.all;
entity memory2_vlg_sample_tst is
    port(
        bcd             : in     vl_logic_vector(3 downto 0);
        sampler_tx      : out    vl_logic
    );
end memory2_vlg_sample_tst;
