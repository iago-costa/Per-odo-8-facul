*** SPICE deck for cell NAND_sim{sch} from library tutorial_4
*** Created on Sun May 15, 2022 22:59:24
*** Last revised on Mon May 16, 2022 00:08:26
*** Written on Mon May 16, 2022 00:08:51 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT tutorial_4__NAND_2 FROM CELL NAND_2{sch}
.SUBCKT tutorial_4__NAND_2 A AnandB B
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 AnandB A net@45 gnd NMOS L=0.6U W=3U
Mnmos@1 AnandB A vdd vdd PMOS L=0.6U W=3U
Mnmos@2 net@45 B gnd gnd NMOS L=0.6U W=3U
Mpmos@0 AnandB B vdd vdd PMOS L=0.6U W=3U
.ENDS tutorial_4__NAND_2

.global gnd vdd

*** TOP LEVEL CELL: NAND_sim{sch}
XNAND_2@1 in out vdd tutorial_4__NAND_2

* Spice Code nodes in cell cell 'NAND_sim{sch}'
vdd vdd 0 dc 5
vin in 0 dc 0 pulse 0 5 10n 1n
cload out 0 250fF
.tran 0 40n
.include c5_models.txt
.END
