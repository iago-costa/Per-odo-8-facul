library verilog;
use verilog.vl_types.all;
entity address_decoder_vlg_vec_tst is
end address_decoder_vlg_vec_tst;
