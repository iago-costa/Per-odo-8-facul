library verilog;
use verilog.vl_types.all;
entity memory4_vlg_vec_tst is
end memory4_vlg_vec_tst;
